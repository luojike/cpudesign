library ieee;
use ieee.std_logic_1164.all;
use work.opcodes.all;
use work.pc.all;

-- Entity main:
-- The core CPU that consists of components defined in different files.
entity main is
    port (
        clk : in std_logic;
        ir : 
    )
end main;