library ieee;
use ieee.numeric_bit.all;

package myprober is
	signal test : unsigned(31 downto 0) := X"00000000";
end package myprober;
